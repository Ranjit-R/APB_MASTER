`define data_width 32
`define addr_width 8
`define strb_width data_width/8

`define no_trans 10

